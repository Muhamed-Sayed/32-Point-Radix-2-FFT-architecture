module FFT_module(X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,X16,X17,X18,X19,X20,X21,X22,X23,
				  X24,X25,X26,X27,X28,X29,X30,X31,
				  	S5_OUT0r_reg,S5_OUT0i_reg,S5_OUT1r_reg,S5_OUT1i_reg,S5_OUT2r_reg,S5_OUT2i_reg,S5_OUT3r_reg,S5_OUT3i_reg,S5_OUT4r_reg,S5_OUT4i_reg,
			S5_OUT5r_reg,S5_OUT5i_reg,S5_OUT6r_reg,S5_OUT6i_reg,S5_OUT7r_reg,S5_OUT7i_reg,S5_OUT8r_reg,S5_OUT8i_reg,S5_OUT9r_reg,S5_OUT9i_reg,
			S5_OUT10r_reg,S5_OUT10i_reg,S5_OUT11r_reg,S5_OUT11i_reg,S5_OUT12r_reg,S5_OUT12i_reg,S5_OUT13r_reg,S5_OUT13i_reg,S5_OUT14r_reg,
			S5_OUT14i_reg,S5_OUT15r_reg,S5_OUT15i_reg,S5_OUT16r_reg,S5_OUT16i_reg,S5_OUT17r_reg,S5_OUT17i_reg,S5_OUT18r_reg,S5_OUT18i_reg,
			S5_OUT19r_reg,S5_OUT19i_reg,S5_OUT20r_reg,S5_OUT20i_reg,S5_OUT21r_reg,S5_OUT21i_reg,S5_OUT22r_reg,S5_OUT22i_reg,S5_OUT23r_reg,
			S5_OUT23i_reg,S5_OUT24r_reg,S5_OUT24i_reg,S5_OUT25r_reg,S5_OUT25i_reg,S5_OUT26r_reg,S5_OUT26i_reg,S5_OUT27r_reg,S5_OUT27i_reg,
			S5_OUT28r_reg,S5_OUT28i_reg,S5_OUT29r_reg,S5_OUT29i_reg,S5_OUT30r_reg,S5_OUT30i_reg,S5_OUT31r_reg,S5_OUT31i_reg,
				  clk,clk_MAC,rst);

input wire clk,clk_MAC,rst;
input wire [7:0] X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,X16,X17,X18,X19,X20,X21,X22,X23,X24,X25,X26,X27,X28,X29,X30,X31;
output wire [15:0]	S5_OUT0r_reg,S5_OUT0i_reg,S5_OUT1r_reg,S5_OUT1i_reg,S5_OUT2r_reg,S5_OUT2i_reg,S5_OUT3r_reg,S5_OUT3i_reg,S5_OUT4r_reg,S5_OUT4i_reg,
			S5_OUT5r_reg,S5_OUT5i_reg,S5_OUT6r_reg,S5_OUT6i_reg,S5_OUT7r_reg,S5_OUT7i_reg,S5_OUT8r_reg,S5_OUT8i_reg,S5_OUT9r_reg,S5_OUT9i_reg,
			S5_OUT10r_reg,S5_OUT10i_reg,S5_OUT11r_reg,S5_OUT11i_reg,S5_OUT12r_reg,S5_OUT12i_reg,S5_OUT13r_reg,S5_OUT13i_reg,S5_OUT14r_reg,
			S5_OUT14i_reg,S5_OUT15r_reg,S5_OUT15i_reg,S5_OUT16r_reg,S5_OUT16i_reg,S5_OUT17r_reg,S5_OUT17i_reg,S5_OUT18r_reg,S5_OUT18i_reg,
			S5_OUT19r_reg,S5_OUT19i_reg,S5_OUT20r_reg,S5_OUT20i_reg,S5_OUT21r_reg,S5_OUT21i_reg,S5_OUT22r_reg,S5_OUT22i_reg,S5_OUT23r_reg,
			S5_OUT23i_reg,S5_OUT24r_reg,S5_OUT24i_reg,S5_OUT25r_reg,S5_OUT25i_reg,S5_OUT26r_reg,S5_OUT26i_reg,S5_OUT27r_reg,S5_OUT27i_reg,
			S5_OUT28r_reg,S5_OUT28i_reg,S5_OUT29r_reg,S5_OUT29i_reg,S5_OUT30r_reg,S5_OUT30i_reg,S5_OUT31r_reg,S5_OUT31i_reg;

wire [15:0] W0r,W0i,W1r,W1i,W2r,W2i,W3r,W3i,W4r,W4i,W5r,W5i,W6r,W6i,W7r,W7i,
		   W8r,W8i,W9r,W9i,W10r,W10i,W11r,W11i,W12r,W12i,W13r,W13i,W14r,W14i,W15r,W15i;

wire [15:0] 	S1_OUT0r,S1_OUT0i,S1_OUT1r,S1_OUT1i,S1_OUT2r,S1_OUT2i,S1_OUT3r,S1_OUT3i,S1_OUT4r,S1_OUT4i,
			S1_OUT5r,S1_OUT5i,S1_OUT6r,S1_OUT6i,S1_OUT7r,S1_OUT7i,S1_OUT8r,S1_OUT8i,S1_OUT9r,S1_OUT9i,
			S1_OUT10r,S1_OUT10i,S1_OUT11r,S1_OUT11i,S1_OUT12r,S1_OUT12i,S1_OUT13r,S1_OUT13i,S1_OUT14r,
			S1_OUT14i,S1_OUT15r,S1_OUT15i,S1_OUT16r,S1_OUT16i,S1_OUT17r,S1_OUT17i,S1_OUT18r,S1_OUT18i,
			S1_OUT19r,S1_OUT19i,S1_OUT20r,S1_OUT20i,S1_OUT21r,S1_OUT21i,S1_OUT22r,S1_OUT22i,S1_OUT23r,
			S1_OUT23i,S1_OUT24r,S1_OUT24i,S1_OUT25r,S1_OUT25i,S1_OUT26r,S1_OUT26i,S1_OUT27r,S1_OUT27i,
			S1_OUT28r,S1_OUT28i,S1_OUT29r,S1_OUT29i,S1_OUT30r,S1_OUT30i,S1_OUT31r,S1_OUT31i,
			S2_OUT0r,S2_OUT0i,S2_OUT1r,S2_OUT1i,S2_OUT2r,S2_OUT2i,S2_OUT3r,S2_OUT3i,S2_OUT4r,S2_OUT4i,
			S2_OUT5r,S2_OUT5i,S2_OUT6r,S2_OUT6i,S2_OUT7r,S2_OUT7i,S2_OUT8r,S2_OUT8i,S2_OUT9r,S2_OUT9i,
			S2_OUT10r,S2_OUT10i,S2_OUT11r,S2_OUT11i,S2_OUT12r,S2_OUT12i,S2_OUT13r,S2_OUT13i,S2_OUT14r,
			S2_OUT14i,S2_OUT15r,S2_OUT15i,S2_OUT16r,S2_OUT16i,S2_OUT17r,S2_OUT17i,S2_OUT18r,S2_OUT18i,
			S2_OUT19r,S2_OUT19i,S2_OUT20r,S2_OUT20i,S2_OUT21r,S2_OUT21i,S2_OUT22r,S2_OUT22i,S2_OUT23r,
			S2_OUT23i,S2_OUT24r,S2_OUT24i,S2_OUT25r,S2_OUT25i,S2_OUT26r,S2_OUT26i,S2_OUT27r,S2_OUT27i,
			S2_OUT28r,S2_OUT28i,S2_OUT29r,S2_OUT29i,S2_OUT30r,S2_OUT30i,S2_OUT31r,S2_OUT31i,
			S3_OUT0r,S3_OUT0i,S3_OUT1r,S3_OUT1i,S3_OUT2r,S3_OUT2i,S3_OUT3r,S3_OUT3i,S3_OUT4r,S3_OUT4i,
			S3_OUT5r,S3_OUT5i,S3_OUT6r,S3_OUT6i,S3_OUT7r,S3_OUT7i,S3_OUT8r,S3_OUT8i,S3_OUT9r,S3_OUT9i,
			S3_OUT10r,S3_OUT10i,S3_OUT11r,S3_OUT11i,S3_OUT12r,S3_OUT12i,S3_OUT13r,S3_OUT13i,S3_OUT14r,
			S3_OUT14i,S3_OUT15r,S3_OUT15i,S3_OUT16r,S3_OUT16i,S3_OUT17r,S3_OUT17i,S3_OUT18r,S3_OUT18i,
			S3_OUT19r,S3_OUT19i,S3_OUT20r,S3_OUT20i,S3_OUT21r,S3_OUT21i,S3_OUT22r,S3_OUT22i,S3_OUT23r,
			S3_OUT23i,S3_OUT24r,S3_OUT24i,S3_OUT25r,S3_OUT25i,S3_OUT26r,S3_OUT26i,S3_OUT27r,S3_OUT27i,
			S3_OUT28r,S3_OUT28i,S3_OUT29r,S3_OUT29i,S3_OUT30r,S3_OUT30i,S3_OUT31r,S3_OUT31i,
			S4_OUT0r,S4_OUT0i,S4_OUT1r,S4_OUT1i,S4_OUT2r,S4_OUT2i,S4_OUT3r,S4_OUT3i,S4_OUT4r,S4_OUT4i,
			S4_OUT5r,S4_OUT5i,S4_OUT6r,S4_OUT6i,S4_OUT7r,S4_OUT7i,S4_OUT8r,S4_OUT8i,S4_OUT9r,S4_OUT9i,
			S4_OUT10r,S4_OUT10i,S4_OUT11r,S4_OUT11i,S4_OUT12r,S4_OUT12i,S4_OUT13r,S4_OUT13i,S4_OUT14r,
			S4_OUT14i,S4_OUT15r,S4_OUT15i,S4_OUT16r,S4_OUT16i,S4_OUT17r,S4_OUT17i,S4_OUT18r,S4_OUT18i,
			S4_OUT19r,S4_OUT19i,S4_OUT20r,S4_OUT20i,S4_OUT21r,S4_OUT21i,S4_OUT22r,S4_OUT22i,S4_OUT23r,
			S4_OUT23i,S4_OUT24r,S4_OUT24i,S4_OUT25r,S4_OUT25i,S4_OUT26r,S4_OUT26i,S4_OUT27r,S4_OUT27i,
			S4_OUT28r,S4_OUT28i,S4_OUT29r,S4_OUT29i,S4_OUT30r,S4_OUT30i,S4_OUT31r,S4_OUT31i,
			S5_OUT0r,S5_OUT0i,S5_OUT1r,S5_OUT1i,S5_OUT2r,S5_OUT2i,S5_OUT3r,S5_OUT3i,S5_OUT4r,S5_OUT4i,S5_OUT5r,S5_OUT5i,
			S5_OUT6r,S5_OUT6i,S5_OUT7r,S5_OUT7i,S5_OUT8r,S5_OUT8i,S5_OUT9r,S5_OUT9i,S5_OUT10r,S5_OUT10i,S5_OUT11r,S5_OUT11i,
			S5_OUT12r,S5_OUT12i,S5_OUT13r,S5_OUT13i,S5_OUT14r,S5_OUT14i,S5_OUT15r,S5_OUT15i,S5_OUT16r,S5_OUT16i,S5_OUT17r,
			S5_OUT17i,S5_OUT18r,S5_OUT18i,S5_OUT19r,S5_OUT19i,S5_OUT20r,S5_OUT20i,S5_OUT21r,S5_OUT21i,S5_OUT22r,S5_OUT22i,
			S5_OUT23r,S5_OUT23i,S5_OUT24r,S5_OUT24i,S5_OUT25r,S5_OUT25i,S5_OUT26r,S5_OUT26i,S5_OUT27r,S5_OUT27i,S5_OUT28r,
			S5_OUT28i,S5_OUT29r,S5_OUT29i,S5_OUT30r,S5_OUT30i,S5_OUT31r,S5_OUT31i,
			S1_OUT0r_reg,S1_OUT0i_reg,S1_OUT1r_reg,S1_OUT1i_reg,S1_OUT2r_reg,S1_OUT2i_reg,S1_OUT3r_reg,S1_OUT3i_reg,S1_OUT4r_reg,S1_OUT4i_reg,
			S1_OUT5r_reg,S1_OUT5i_reg,S1_OUT6r_reg,S1_OUT6i_reg,S1_OUT7r_reg,S1_OUT7i_reg,S1_OUT8r_reg,S1_OUT8i_reg,S1_OUT9r_reg,S1_OUT9i_reg,
			S1_OUT10r_reg,S1_OUT10i_reg,S1_OUT11r_reg,S1_OUT11i_reg,S1_OUT12r_reg,S1_OUT12i_reg,S1_OUT13r_reg,S1_OUT13i_reg,S1_OUT14r_reg,
			S1_OUT14i_reg,S1_OUT15r_reg,S1_OUT15i_reg,S1_OUT16r_reg,S1_OUT16i_reg,S1_OUT17r_reg,S1_OUT17i_reg,S1_OUT18r_reg,S1_OUT18i_reg,
			S1_OUT19r_reg,S1_OUT19i_reg,S1_OUT20r_reg,S1_OUT20i_reg,S1_OUT21r_reg,S1_OUT21i_reg,S1_OUT22r_reg,S1_OUT22i_reg,S1_OUT23r_reg,
			S1_OUT23i_reg,S1_OUT24r_reg,S1_OUT24i_reg,S1_OUT25r_reg,S1_OUT25i_reg,S1_OUT26r_reg,S1_OUT26i_reg,S1_OUT27r_reg,S1_OUT27i_reg,
			S1_OUT28r_reg,S1_OUT28i_reg,S1_OUT29r_reg,S1_OUT29i_reg,S1_OUT30r_reg,S1_OUT30i_reg,S1_OUT31r_reg,S1_OUT31i_reg,
			S2_OUT0r_reg,S2_OUT0i_reg,S2_OUT1r_reg,S2_OUT1i_reg,S2_OUT2r_reg,S2_OUT2i_reg,S2_OUT3r_reg,S2_OUT3i_reg,S2_OUT4r_reg,S2_OUT4i_reg,
			S2_OUT5r_reg,S2_OUT5i_reg,S2_OUT6r_reg,S2_OUT6i_reg,S2_OUT7r_reg,S2_OUT7i_reg,S2_OUT8r_reg,S2_OUT8i_reg,S2_OUT9r_reg,S2_OUT9i_reg,
			S2_OUT10r_reg,S2_OUT10i_reg,S2_OUT11r_reg,S2_OUT11i_reg,S2_OUT12r_reg,S2_OUT12i_reg,S2_OUT13r_reg,S2_OUT13i_reg,S2_OUT14r_reg,
			S2_OUT14i_reg,S2_OUT15r_reg,S2_OUT15i_reg,S2_OUT16r_reg,S2_OUT16i_reg,S2_OUT17r_reg,S2_OUT17i_reg,S2_OUT18r_reg,S2_OUT18i_reg,
			S2_OUT19r_reg,S2_OUT19i_reg,S2_OUT20r_reg,S2_OUT20i_reg,S2_OUT21r_reg,S2_OUT21i_reg,S2_OUT22r_reg,S2_OUT22i_reg,S2_OUT23r_reg,
			S2_OUT23i_reg,S2_OUT24r_reg,S2_OUT24i_reg,S2_OUT25r_reg,S2_OUT25i_reg,S2_OUT26r_reg,S2_OUT26i_reg,S2_OUT27r_reg,S2_OUT27i_reg,
			S2_OUT28r_reg,S2_OUT28i_reg,S2_OUT29r_reg,S2_OUT29i_reg,S2_OUT30r_reg,S2_OUT30i_reg,S2_OUT31r_reg,S2_OUT31i_reg,
			S3_OUT0r_reg,S3_OUT0i_reg,S3_OUT1r_reg,S3_OUT1i_reg,S3_OUT2r_reg,S3_OUT2i_reg,S3_OUT3r_reg,S3_OUT3i_reg,S3_OUT4r_reg,S3_OUT4i_reg,
			S3_OUT5r_reg,S3_OUT5i_reg,S3_OUT6r_reg,S3_OUT6i_reg,S3_OUT7r_reg,S3_OUT7i_reg,S3_OUT8r_reg,S3_OUT8i_reg,S3_OUT9r_reg,S3_OUT9i_reg,
			S3_OUT10r_reg,S3_OUT10i_reg,S3_OUT11r_reg,S3_OUT11i_reg,S3_OUT12r_reg,S3_OUT12i_reg,S3_OUT13r_reg,S3_OUT13i_reg,S3_OUT14r_reg,
			S3_OUT14i_reg,S3_OUT15r_reg,S3_OUT15i_reg,S3_OUT16r_reg,S3_OUT16i_reg,S3_OUT17r_reg,S3_OUT17i_reg,S3_OUT18r_reg,S3_OUT18i_reg,
			S3_OUT19r_reg,S3_OUT19i_reg,S3_OUT20r_reg,S3_OUT20i_reg,S3_OUT21r_reg,S3_OUT21i_reg,S3_OUT22r_reg,S3_OUT22i_reg,S3_OUT23r_reg,
			S3_OUT23i_reg,S3_OUT24r_reg,S3_OUT24i_reg,S3_OUT25r_reg,S3_OUT25i_reg,S3_OUT26r_reg,S3_OUT26i_reg,S3_OUT27r_reg,S3_OUT27i_reg,
			S3_OUT28r_reg,S3_OUT28i_reg,S3_OUT29r_reg,S3_OUT29i_reg,S3_OUT30r_reg,S3_OUT30i_reg,S3_OUT31r_reg,S3_OUT31i_reg,
			S4_OUT0r_reg,S4_OUT0i_reg,S4_OUT1r_reg,S4_OUT1i_reg,S4_OUT2r_reg,S4_OUT2i_reg,S4_OUT3r_reg,S4_OUT3i_reg,S4_OUT4r_reg,S4_OUT4i_reg,
			S4_OUT5r_reg,S4_OUT5i_reg,S4_OUT6r_reg,S4_OUT6i_reg,S4_OUT7r_reg,S4_OUT7i_reg,S4_OUT8r_reg,S4_OUT8i_reg,S4_OUT9r_reg,S4_OUT9i_reg,
			S4_OUT10r_reg,S4_OUT10i_reg,S4_OUT11r_reg,S4_OUT11i_reg,S4_OUT12r_reg,S4_OUT12i_reg,S4_OUT13r_reg,S4_OUT13i_reg,S4_OUT14r_reg,
			S4_OUT14i_reg,S4_OUT15r_reg,S4_OUT15i_reg,S4_OUT16r_reg,S4_OUT16i_reg,S4_OUT17r_reg,S4_OUT17i_reg,S4_OUT18r_reg,S4_OUT18i_reg,
			S4_OUT19r_reg,S4_OUT19i_reg,S4_OUT20r_reg,S4_OUT20i_reg,S4_OUT21r_reg,S4_OUT21i_reg,S4_OUT22r_reg,S4_OUT22i_reg,S4_OUT23r_reg,
			S4_OUT23i_reg,S4_OUT24r_reg,S4_OUT24i_reg,S4_OUT25r_reg,S4_OUT25i_reg,S4_OUT26r_reg,S4_OUT26i_reg,S4_OUT27r_reg,S4_OUT27i_reg,
			S4_OUT28r_reg,S4_OUT28i_reg,S4_OUT29r_reg,S4_OUT29i_reg,S4_OUT30r_reg,S4_OUT30i_reg,S4_OUT31r_reg,S4_OUT31i_reg;
			
wire [2:0] count,count_reg;
wire flag;

counter counter(clk_MAC,count,rst);
reg_count reg_count(count,count_reg,clk_MAC,flag,rst);
			  
memory_W memory_W(W0r,W1r,W2r,W3r,W4r,W5r,W6r,W7r,W8r,W9r,W10r,W11r,W12r,W13r,W14r,W15r,
				  W0i,W1i,W2i,W3i,W4i,W5i,W6i,W7i,W8i,W9i,W10i,W11i,W12i,W13i,W14i,W15i);

stage1 s1(X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,X16,X17,X18,X19,X20,X21,X22,X23,X24,X25,X26,X27,X28,X29,X30,X31,
		  W0r,W0i,
		  S1_OUT0r,S1_OUT0i,S1_OUT1r,S1_OUT1i,S1_OUT2r,S1_OUT2i,S1_OUT3r,S1_OUT3i,S1_OUT4r,S1_OUT4i,S1_OUT5r,S1_OUT5i,S1_OUT6r,S1_OUT6i,
	      S1_OUT7r,S1_OUT7i,S1_OUT8r,S1_OUT8i,S1_OUT9r,S1_OUT9i,S1_OUT10r,S1_OUT10i,S1_OUT11r,S1_OUT11i,S1_OUT12r,S1_OUT12i,S1_OUT13r,S1_OUT13i,
		  S1_OUT14r,S1_OUT14i,S1_OUT15r,S1_OUT15i,S1_OUT16r,S1_OUT16i,S1_OUT17r,S1_OUT17i,S1_OUT18r,S1_OUT18i,S1_OUT19r,S1_OUT19i,S1_OUT20r,
		  S1_OUT20i,S1_OUT21r,S1_OUT21i,S1_OUT22r,S1_OUT22i,S1_OUT23r,S1_OUT23i,S1_OUT24r,S1_OUT24i,S1_OUT25r,S1_OUT25i,S1_OUT26r,S1_OUT26i,
		  S1_OUT27r,S1_OUT27i,S1_OUT28r,S1_OUT28i,S1_OUT29r,S1_OUT29i,S1_OUT30r,S1_OUT30i,S1_OUT31r,S1_OUT31i,clk_MAC,rst,count_reg,count,flag);			
			 
Register #(.size(16)) Register_S1_0(S1_OUT0r,S1_OUT0i,S1_OUT0r_reg,S1_OUT0i_reg,clk,rst);
Register #(.size(16)) Register_S1_1(S1_OUT1r,S1_OUT1i,S1_OUT1r_reg,S1_OUT1i_reg,clk,rst);
Register #(.size(16)) Register_S1_2(S1_OUT2r,S1_OUT2i,S1_OUT2r_reg,S1_OUT2i_reg,clk,rst);
Register #(.size(16)) Register_S1_3(S1_OUT3r,S1_OUT3i,S1_OUT3r_reg,S1_OUT3i_reg,clk,rst);
Register #(.size(16)) Register_S1_4(S1_OUT4r,S1_OUT4i,S1_OUT4r_reg,S1_OUT4i_reg,clk,rst);
Register #(.size(16)) Register_S1_5(S1_OUT5r,S1_OUT5i,S1_OUT5r_reg,S1_OUT5i_reg,clk,rst);
Register #(.size(16)) Register_S1_6(S1_OUT6r,S1_OUT6i,S1_OUT6r_reg,S1_OUT6i_reg,clk,rst);
Register #(.size(16)) Register_S1_7(S1_OUT7r,S1_OUT7i,S1_OUT7r_reg,S1_OUT7i_reg,clk,rst);
Register #(.size(16)) Register_S1_8(S1_OUT8r,S1_OUT8i,S1_OUT8r_reg,S1_OUT8i_reg,clk,rst);
Register #(.size(16)) Register_S1_9(S1_OUT9r,S1_OUT9i,S1_OUT9r_reg,S1_OUT9i_reg,clk,rst);
Register #(.size(16)) Register_S1_10(S1_OUT10r,S1_OUT10i,S1_OUT10r_reg,S1_OUT10i_reg,clk,rst);
Register #(.size(16)) Register_S1_11(S1_OUT11r,S1_OUT11i,S1_OUT11r_reg,S1_OUT11i_reg,clk,rst);
Register #(.size(16)) Register_S1_12(S1_OUT12r,S1_OUT12i,S1_OUT12r_reg,S1_OUT12i_reg,clk,rst);
Register #(.size(16)) Register_S1_13(S1_OUT13r,S1_OUT13i,S1_OUT13r_reg,S1_OUT13i_reg,clk,rst);
Register #(.size(16)) Register_S1_14(S1_OUT14r,S1_OUT14i,S1_OUT14r_reg,S1_OUT14i_reg,clk,rst);
Register #(.size(16)) Register_S1_15(S1_OUT15r,S1_OUT15i,S1_OUT15r_reg,S1_OUT15i_reg,clk,rst);
Register #(.size(16)) Register_S1_16(S1_OUT16r,S1_OUT16i,S1_OUT16r_reg,S1_OUT16i_reg,clk,rst);
Register #(.size(16)) Register_S1_17(S1_OUT17r,S1_OUT17i,S1_OUT17r_reg,S1_OUT17i_reg,clk,rst);
Register #(.size(16)) Register_S1_18(S1_OUT18r,S1_OUT18i,S1_OUT18r_reg,S1_OUT18i_reg,clk,rst);
Register #(.size(16)) Register_S1_19(S1_OUT19r,S1_OUT19i,S1_OUT19r_reg,S1_OUT19i_reg,clk,rst);
Register #(.size(16)) Register_S1_20(S1_OUT20r,S1_OUT20i,S1_OUT20r_reg,S1_OUT20i_reg,clk,rst);
Register #(.size(16)) Register_S1_21(S1_OUT21r,S1_OUT21i,S1_OUT21r_reg,S1_OUT21i_reg,clk,rst);
Register #(.size(16)) Register_S1_22(S1_OUT22r,S1_OUT22i,S1_OUT22r_reg,S1_OUT22i_reg,clk,rst);
Register #(.size(16)) Register_S1_23(S1_OUT23r,S1_OUT23i,S1_OUT23r_reg,S1_OUT23i_reg,clk,rst);
Register #(.size(16)) Register_S1_24(S1_OUT24r,S1_OUT24i,S1_OUT24r_reg,S1_OUT24i_reg,clk,rst);
Register #(.size(16)) Register_S1_25(S1_OUT25r,S1_OUT25i,S1_OUT25r_reg,S1_OUT25i_reg,clk,rst);
Register #(.size(16)) Register_S1_26(S1_OUT26r,S1_OUT26i,S1_OUT26r_reg,S1_OUT26i_reg,clk,rst);
Register #(.size(16)) Register_S1_27(S1_OUT27r,S1_OUT27i,S1_OUT27r_reg,S1_OUT27i_reg,clk,rst);
Register #(.size(16)) Register_S1_28(S1_OUT28r,S1_OUT28i,S1_OUT28r_reg,S1_OUT28i_reg,clk,rst);
Register #(.size(16)) Register_S1_29(S1_OUT29r,S1_OUT29i,S1_OUT29r_reg,S1_OUT29i_reg,clk,rst);
Register #(.size(16)) Register_S1_30(S1_OUT30r,S1_OUT30i,S1_OUT30r_reg,S1_OUT30i_reg,clk,rst);
Register #(.size(16)) Register_S1_31(S1_OUT31r,S1_OUT31i,S1_OUT31r_reg,S1_OUT31i_reg,clk,rst);

stage2 S2(S1_OUT0r_reg,S1_OUT0i_reg,S1_OUT1r_reg,S1_OUT1i_reg,S1_OUT2r_reg,S1_OUT2i_reg,S1_OUT3r_reg,S1_OUT3i_reg,
		  S1_OUT4r_reg,S1_OUT4i_reg,S1_OUT5r_reg,S1_OUT5i_reg,S1_OUT6r_reg,S1_OUT6i_reg,S1_OUT7r_reg,S1_OUT7i_reg,
		  S1_OUT8r_reg,S1_OUT8i_reg,S1_OUT9r_reg,S1_OUT9i_reg,S1_OUT10r_reg,S1_OUT10i_reg,S1_OUT11r_reg,S1_OUT11i_reg,
		  S1_OUT12r_reg,S1_OUT12i_reg,S1_OUT13r_reg,S1_OUT13i_reg,S1_OUT14r_reg,S1_OUT14i_reg,S1_OUT15r_reg,S1_OUT15i_reg,
		  S1_OUT16r_reg,S1_OUT16i_reg,S1_OUT17r_reg,S1_OUT17i_reg,S1_OUT18r_reg,S1_OUT18i_reg,S1_OUT19r_reg,S1_OUT19i_reg,
		  S1_OUT20r_reg,S1_OUT20i_reg,S1_OUT21r_reg,S1_OUT21i_reg,S1_OUT22r_reg,S1_OUT22i_reg,S1_OUT23r_reg,S1_OUT23i_reg,
		  S1_OUT24r_reg,S1_OUT24i_reg,S1_OUT25r_reg,S1_OUT25i_reg,S1_OUT26r_reg,S1_OUT26i_reg,S1_OUT27r_reg,S1_OUT27i_reg,
		  S1_OUT28r_reg,S1_OUT28i_reg,S1_OUT29r_reg,S1_OUT29i_reg,S1_OUT30r_reg,S1_OUT30i_reg,S1_OUT31r_reg,S1_OUT31i_reg,
		  W0r,W0i,W8r,W8i,
		  S2_OUT0r,S2_OUT0i,S2_OUT1r,S2_OUT1i,S2_OUT2r,S2_OUT2i,S2_OUT3r,S2_OUT3i,S2_OUT4r,S2_OUT4i,S2_OUT5r,S2_OUT5i,
		  S2_OUT6r,S2_OUT6i,S2_OUT7r,S2_OUT7i,S2_OUT8r,S2_OUT8i,S2_OUT9r,S2_OUT9i,S2_OUT10r,S2_OUT10i,S2_OUT11r,S2_OUT11i,
		  S2_OUT12r,S2_OUT12i,S2_OUT13r,S2_OUT13i,S2_OUT14r,S2_OUT14i,S2_OUT15r,S2_OUT15i,S2_OUT16r,S2_OUT16i,S2_OUT17r,
		  S2_OUT17i,S2_OUT18r,S2_OUT18i,S2_OUT19r,S2_OUT19i,S2_OUT20r,S2_OUT20i,S2_OUT21r,S2_OUT21i,S2_OUT22r,S2_OUT22i,
		  S2_OUT23r,S2_OUT23i,S2_OUT24r,S2_OUT24i,S2_OUT25r,S2_OUT25i,S2_OUT26r,S2_OUT26i,S2_OUT27r,S2_OUT27i,S2_OUT28r,
		  S2_OUT28i,S2_OUT29r,S2_OUT29i,S2_OUT30r,S2_OUT30i,S2_OUT31r,S2_OUT31i,
		  clk_MAC,rst,count_reg,count,flag);	
			 
Register #(.size(16)) Register_S2_0(S2_OUT0r,S2_OUT0i,S2_OUT0r_reg,S2_OUT0i_reg,clk,rst);
Register #(.size(16)) Register_S2_1(S2_OUT1r,S2_OUT1i,S2_OUT1r_reg,S2_OUT1i_reg,clk,rst);
Register #(.size(16)) Register_S2_2(S2_OUT2r,S2_OUT2i,S2_OUT2r_reg,S2_OUT2i_reg,clk,rst);
Register #(.size(16)) Register_S2_3(S2_OUT3r,S2_OUT3i,S2_OUT3r_reg,S2_OUT3i_reg,clk,rst);
Register #(.size(16)) Register_S2_4(S2_OUT4r,S2_OUT4i,S2_OUT4r_reg,S2_OUT4i_reg,clk,rst);
Register #(.size(16)) Register_S2_5(S2_OUT5r,S2_OUT5i,S2_OUT5r_reg,S2_OUT5i_reg,clk,rst);
Register #(.size(16)) Register_S2_6(S2_OUT6r,S2_OUT6i,S2_OUT6r_reg,S2_OUT6i_reg,clk,rst);
Register #(.size(16)) Register_S2_7(S2_OUT7r,S2_OUT7i,S2_OUT7r_reg,S2_OUT7i_reg,clk,rst);
Register #(.size(16)) Register_S2_8(S2_OUT8r,S2_OUT8i,S2_OUT8r_reg,S2_OUT8i_reg,clk,rst);
Register #(.size(16)) Register_S2_9(S2_OUT9r,S2_OUT9i,S2_OUT9r_reg,S2_OUT9i_reg,clk,rst);
Register #(.size(16)) Register_S2_10(S2_OUT10r,S2_OUT10i,S2_OUT10r_reg,S2_OUT10i_reg,clk,rst);
Register #(.size(16)) Register_S2_11(S2_OUT11r,S2_OUT11i,S2_OUT11r_reg,S2_OUT11i_reg,clk,rst);
Register #(.size(16)) Register_S2_12(S2_OUT12r,S2_OUT12i,S2_OUT12r_reg,S2_OUT12i_reg,clk,rst);
Register #(.size(16)) Register_S2_13(S2_OUT13r,S2_OUT13i,S2_OUT13r_reg,S2_OUT13i_reg,clk,rst);
Register #(.size(16)) Register_S2_14(S2_OUT14r,S2_OUT14i,S2_OUT14r_reg,S2_OUT14i_reg,clk,rst);
Register #(.size(16)) Register_S2_15(S2_OUT15r,S2_OUT15i,S2_OUT15r_reg,S2_OUT15i_reg,clk,rst);
Register #(.size(16)) Register_S2_16(S2_OUT16r,S2_OUT16i,S2_OUT16r_reg,S2_OUT16i_reg,clk,rst);
Register #(.size(16)) Register_S2_17(S2_OUT17r,S2_OUT17i,S2_OUT17r_reg,S2_OUT17i_reg,clk,rst);
Register #(.size(16)) Register_S2_18(S2_OUT18r,S2_OUT18i,S2_OUT18r_reg,S2_OUT18i_reg,clk,rst);
Register #(.size(16)) Register_S2_19(S2_OUT19r,S2_OUT19i,S2_OUT19r_reg,S2_OUT19i_reg,clk,rst);
Register #(.size(16)) Register_S2_20(S2_OUT20r,S2_OUT20i,S2_OUT20r_reg,S2_OUT20i_reg,clk,rst);
Register #(.size(16)) Register_S2_21(S2_OUT21r,S2_OUT21i,S2_OUT21r_reg,S2_OUT21i_reg,clk,rst);
Register #(.size(16)) Register_S2_22(S2_OUT22r,S2_OUT22i,S2_OUT22r_reg,S2_OUT22i_reg,clk,rst);
Register #(.size(16)) Register_S2_23(S2_OUT23r,S2_OUT23i,S2_OUT23r_reg,S2_OUT23i_reg,clk,rst);
Register #(.size(16)) Register_S2_24(S2_OUT24r,S2_OUT24i,S2_OUT24r_reg,S2_OUT24i_reg,clk,rst);
Register #(.size(16)) Register_S2_25(S2_OUT25r,S2_OUT25i,S2_OUT25r_reg,S2_OUT25i_reg,clk,rst);
Register #(.size(16)) Register_S2_26(S2_OUT26r,S2_OUT26i,S2_OUT26r_reg,S2_OUT26i_reg,clk,rst);
Register #(.size(16)) Register_S2_27(S2_OUT27r,S2_OUT27i,S2_OUT27r_reg,S2_OUT27i_reg,clk,rst);
Register #(.size(16)) Register_S2_28(S2_OUT28r,S2_OUT28i,S2_OUT28r_reg,S2_OUT28i_reg,clk,rst);
Register #(.size(16)) Register_S2_29(S2_OUT29r,S2_OUT29i,S2_OUT29r_reg,S2_OUT29i_reg,clk,rst);
Register #(.size(16)) Register_S2_30(S2_OUT30r,S2_OUT30i,S2_OUT30r_reg,S2_OUT30i_reg,clk,rst);
Register #(.size(16)) Register_S2_31(S2_OUT31r,S2_OUT31i,S2_OUT31r_reg,S2_OUT31i_reg,clk,rst);

stage3 S3(S2_OUT0r_reg,S2_OUT0i_reg,S2_OUT1r_reg,S2_OUT1i_reg,S2_OUT2r_reg,S2_OUT2i_reg,S2_OUT3r_reg,S2_OUT3i_reg,
		  S2_OUT4r_reg,S2_OUT4i_reg,S2_OUT5r_reg,S2_OUT5i_reg,S2_OUT6r_reg,S2_OUT6i_reg,S2_OUT7r_reg,S2_OUT7i_reg,
		  S2_OUT8r_reg,S2_OUT8i_reg,S2_OUT9r_reg,S2_OUT9i_reg,S2_OUT10r_reg,S2_OUT10i_reg,S2_OUT11r_reg,S2_OUT11i_reg,
		  S2_OUT12r_reg,S2_OUT12i_reg,S2_OUT13r_reg,S2_OUT13i_reg,S2_OUT14r_reg,S2_OUT14i_reg,S2_OUT15r_reg,S2_OUT15i_reg,
		  S2_OUT16r_reg,S2_OUT16i_reg,S2_OUT17r_reg,S2_OUT17i_reg,S2_OUT18r_reg,S2_OUT18i_reg,S2_OUT19r_reg,S2_OUT19i_reg,
		  S2_OUT20r_reg,S2_OUT20i_reg,S2_OUT21r_reg,S2_OUT21i_reg,S2_OUT22r_reg,S2_OUT22i_reg,S2_OUT23r_reg,S2_OUT23i_reg,
		  S2_OUT24r_reg,S2_OUT24i_reg,S2_OUT25r_reg,S2_OUT25i_reg,S2_OUT26r_reg,S2_OUT26i_reg,S2_OUT27r_reg,S2_OUT27i_reg,
		  S2_OUT28r_reg,S2_OUT28i_reg,S2_OUT29r_reg,S2_OUT29i_reg,S2_OUT30r_reg,S2_OUT30i_reg,S2_OUT31r_reg,S2_OUT31i_reg,
		  W0r,W0i,W4r,W4i,W8r,W8i,W12r,W12i,
		  S3_OUT0r,S3_OUT0i,S3_OUT1r,S3_OUT1i,S3_OUT2r,S3_OUT2i,S3_OUT3r,S3_OUT3i,S3_OUT4r,S3_OUT4i,S3_OUT5r,S3_OUT5i,
		  S3_OUT6r,S3_OUT6i,S3_OUT7r,S3_OUT7i,S3_OUT8r,S3_OUT8i,S3_OUT9r,S3_OUT9i,S3_OUT10r,S3_OUT10i,S3_OUT11r,S3_OUT11i,
		  S3_OUT12r,S3_OUT12i,S3_OUT13r,S3_OUT13i,S3_OUT14r,S3_OUT14i,S3_OUT15r,S3_OUT15i,S3_OUT16r,S3_OUT16i,S3_OUT17r,
		  S3_OUT17i,S3_OUT18r,S3_OUT18i,S3_OUT19r,S3_OUT19i,S3_OUT20r,S3_OUT20i,S3_OUT21r,S3_OUT21i,S3_OUT22r,S3_OUT22i,
		  S3_OUT23r,S3_OUT23i,S3_OUT24r,S3_OUT24i,S3_OUT25r,S3_OUT25i,S3_OUT26r,S3_OUT26i,S3_OUT27r,S3_OUT27i,S3_OUT28r,
		  S3_OUT28i,S3_OUT29r,S3_OUT29i,S3_OUT30r,S3_OUT30i,S3_OUT31r,S3_OUT31i,
		  clk_MAC,rst,count_reg,count,flag);	

Register #(.size(16)) Register_S3_0(S3_OUT0r,S3_OUT0i,S3_OUT0r_reg,S3_OUT0i_reg,clk,rst);
Register #(.size(16)) Register_S3_1(S3_OUT1r,S3_OUT1i,S3_OUT1r_reg,S3_OUT1i_reg,clk,rst);
Register #(.size(16)) Register_S3_2(S3_OUT2r,S3_OUT2i,S3_OUT2r_reg,S3_OUT2i_reg,clk,rst);
Register #(.size(16)) Register_S3_3(S3_OUT3r,S3_OUT3i,S3_OUT3r_reg,S3_OUT3i_reg,clk,rst);
Register #(.size(16)) Register_S3_4(S3_OUT4r,S3_OUT4i,S3_OUT4r_reg,S3_OUT4i_reg,clk,rst);
Register #(.size(16)) Register_S3_5(S3_OUT5r,S3_OUT5i,S3_OUT5r_reg,S3_OUT5i_reg,clk,rst);
Register #(.size(16)) Register_S3_6(S3_OUT6r,S3_OUT6i,S3_OUT6r_reg,S3_OUT6i_reg,clk,rst);
Register #(.size(16)) Register_S3_7(S3_OUT7r,S3_OUT7i,S3_OUT7r_reg,S3_OUT7i_reg,clk,rst);
Register #(.size(16)) Register_S3_8(S3_OUT8r,S3_OUT8i,S3_OUT8r_reg,S3_OUT8i_reg,clk,rst);
Register #(.size(16)) Register_S3_9(S3_OUT9r,S3_OUT9i,S3_OUT9r_reg,S3_OUT9i_reg,clk,rst);
Register #(.size(16)) Register_S3_10(S3_OUT10r,S3_OUT10i,S3_OUT10r_reg,S3_OUT10i_reg,clk,rst);
Register #(.size(16)) Register_S3_11(S3_OUT11r,S3_OUT11i,S3_OUT11r_reg,S3_OUT11i_reg,clk,rst);
Register #(.size(16)) Register_S3_12(S3_OUT12r,S3_OUT12i,S3_OUT12r_reg,S3_OUT12i_reg,clk,rst);
Register #(.size(16)) Register_S3_13(S3_OUT13r,S3_OUT13i,S3_OUT13r_reg,S3_OUT13i_reg,clk,rst);
Register #(.size(16)) Register_S3_14(S3_OUT14r,S3_OUT14i,S3_OUT14r_reg,S3_OUT14i_reg,clk,rst);
Register #(.size(16)) Register_S3_15(S3_OUT15r,S3_OUT15i,S3_OUT15r_reg,S3_OUT15i_reg,clk,rst);
Register #(.size(16)) Register_S3_16(S3_OUT16r,S3_OUT16i,S3_OUT16r_reg,S3_OUT16i_reg,clk,rst);
Register #(.size(16)) Register_S3_17(S3_OUT17r,S3_OUT17i,S3_OUT17r_reg,S3_OUT17i_reg,clk,rst);
Register #(.size(16)) Register_S3_18(S3_OUT18r,S3_OUT18i,S3_OUT18r_reg,S3_OUT18i_reg,clk,rst);
Register #(.size(16)) Register_S3_19(S3_OUT19r,S3_OUT19i,S3_OUT19r_reg,S3_OUT19i_reg,clk,rst);
Register #(.size(16)) Register_S3_20(S3_OUT20r,S3_OUT20i,S3_OUT20r_reg,S3_OUT20i_reg,clk,rst);
Register #(.size(16)) Register_S3_21(S3_OUT21r,S3_OUT21i,S3_OUT21r_reg,S3_OUT21i_reg,clk,rst);
Register #(.size(16)) Register_S3_22(S3_OUT22r,S3_OUT22i,S3_OUT22r_reg,S3_OUT22i_reg,clk,rst);
Register #(.size(16)) Register_S3_23(S3_OUT23r,S3_OUT23i,S3_OUT23r_reg,S3_OUT23i_reg,clk,rst);
Register #(.size(16)) Register_S3_24(S3_OUT24r,S3_OUT24i,S3_OUT24r_reg,S3_OUT24i_reg,clk,rst);
Register #(.size(16)) Register_S3_25(S3_OUT25r,S3_OUT25i,S3_OUT25r_reg,S3_OUT25i_reg,clk,rst);
Register #(.size(16)) Register_S3_26(S3_OUT26r,S3_OUT26i,S3_OUT26r_reg,S3_OUT26i_reg,clk,rst);
Register #(.size(16)) Register_S3_27(S3_OUT27r,S3_OUT27i,S3_OUT27r_reg,S3_OUT27i_reg,clk,rst);
Register #(.size(16)) Register_S3_28(S3_OUT28r,S3_OUT28i,S3_OUT28r_reg,S3_OUT28i_reg,clk,rst);
Register #(.size(16)) Register_S3_29(S3_OUT29r,S3_OUT29i,S3_OUT29r_reg,S3_OUT29i_reg,clk,rst);
Register #(.size(16)) Register_S3_30(S3_OUT30r,S3_OUT30i,S3_OUT30r_reg,S3_OUT30i_reg,clk,rst);
Register #(.size(16)) Register_S3_31(S3_OUT31r,S3_OUT31i,S3_OUT31r_reg,S3_OUT31i_reg,clk,rst);	

stage4 S4(S3_OUT0r_reg,S3_OUT0i_reg,S3_OUT1r_reg,S3_OUT1i_reg,S3_OUT2r_reg,S3_OUT2i_reg,S3_OUT3r_reg,S3_OUT3i_reg,
		  S3_OUT4r_reg,S3_OUT4i_reg,S3_OUT5r_reg,S3_OUT5i_reg,S3_OUT6r_reg,S3_OUT6i_reg,S3_OUT7r_reg,S3_OUT7i_reg,
		  S3_OUT8r_reg,S3_OUT8i_reg,S3_OUT9r_reg,S3_OUT9i_reg,S3_OUT10r_reg,S3_OUT10i_reg,S3_OUT11r_reg,S3_OUT11i_reg,
		  S3_OUT12r_reg,S3_OUT12i_reg,S3_OUT13r_reg,S3_OUT13i_reg,S3_OUT14r_reg,S3_OUT14i_reg,S3_OUT15r_reg,S3_OUT15i_reg,
		  S3_OUT16r_reg,S3_OUT16i_reg,S3_OUT17r_reg,S3_OUT17i_reg,S3_OUT18r_reg,S3_OUT18i_reg,S3_OUT19r_reg,S3_OUT19i_reg,
		  S3_OUT20r_reg,S3_OUT20i_reg,S3_OUT21r_reg,S3_OUT21i_reg,S3_OUT22r_reg,S3_OUT22i_reg,S3_OUT23r_reg,S3_OUT23i_reg,
		  S3_OUT24r_reg,S3_OUT24i_reg,S3_OUT25r_reg,S3_OUT25i_reg,S3_OUT26r_reg,S3_OUT26i_reg,S3_OUT27r_reg,S3_OUT27i_reg,
		  S3_OUT28r_reg,S3_OUT28i_reg,S3_OUT29r_reg,S3_OUT29i_reg,S3_OUT30r_reg,S3_OUT30i_reg,S3_OUT31r_reg,S3_OUT31i_reg,
		  W0r,W0i,W2r,W2i,W4r,W4i,W6r,W6i,W8r,W8i,W10r,W10i,W12r,W12i,W14r,W14i,
		  S4_OUT0r,S4_OUT0i,S4_OUT1r,S4_OUT1i,S4_OUT2r,S4_OUT2i,S4_OUT3r,S4_OUT3i,S4_OUT4r,S4_OUT4i,S4_OUT5r,S4_OUT5i,
		  S4_OUT6r,S4_OUT6i,S4_OUT7r,S4_OUT7i,S4_OUT8r,S4_OUT8i,S4_OUT9r,S4_OUT9i,S4_OUT10r,S4_OUT10i,S4_OUT11r,S4_OUT11i,
		  S4_OUT12r,S4_OUT12i,S4_OUT13r,S4_OUT13i,S4_OUT14r,S4_OUT14i,S4_OUT15r,S4_OUT15i,S4_OUT16r,S4_OUT16i,S4_OUT17r,
		  S4_OUT17i,S4_OUT18r,S4_OUT18i,S4_OUT19r,S4_OUT19i,S4_OUT20r,S4_OUT20i,S4_OUT21r,S4_OUT21i,S4_OUT22r,S4_OUT22i,
		  S4_OUT23r,S4_OUT23i,S4_OUT24r,S4_OUT24i,S4_OUT25r,S4_OUT25i,S4_OUT26r,S4_OUT26i,S4_OUT27r,S4_OUT27i,S4_OUT28r,
		  S4_OUT28i,S4_OUT29r,S4_OUT29i,S4_OUT30r,S4_OUT30i,S4_OUT31r,S4_OUT31i,
		  clk_MAC,rst,count_reg,count,flag);	

Register #(.size(16)) Register_S4_0(S4_OUT0r,S4_OUT0i,S4_OUT0r_reg,S4_OUT0i_reg,clk,rst);
Register #(.size(16)) Register_S4_1(S4_OUT1r,S4_OUT1i,S4_OUT1r_reg,S4_OUT1i_reg,clk,rst);
Register #(.size(16)) Register_S4_2(S4_OUT2r,S4_OUT2i,S4_OUT2r_reg,S4_OUT2i_reg,clk,rst);
Register #(.size(16)) Register_S4_3(S4_OUT3r,S4_OUT3i,S4_OUT3r_reg,S4_OUT3i_reg,clk,rst);
Register #(.size(16)) Register_S4_4(S4_OUT4r,S4_OUT4i,S4_OUT4r_reg,S4_OUT4i_reg,clk,rst);
Register #(.size(16)) Register_S4_5(S4_OUT5r,S4_OUT5i,S4_OUT5r_reg,S4_OUT5i_reg,clk,rst);
Register #(.size(16)) Register_S4_6(S4_OUT6r,S4_OUT6i,S4_OUT6r_reg,S4_OUT6i_reg,clk,rst);
Register #(.size(16)) Register_S4_7(S4_OUT7r,S4_OUT7i,S4_OUT7r_reg,S4_OUT7i_reg,clk,rst);
Register #(.size(16)) Register_S4_8(S4_OUT8r,S4_OUT8i,S4_OUT8r_reg,S4_OUT8i_reg,clk,rst);
Register #(.size(16)) Register_S4_9(S4_OUT9r,S4_OUT9i,S4_OUT9r_reg,S4_OUT9i_reg,clk,rst);
Register #(.size(16)) Register_S4_10(S4_OUT10r,S4_OUT10i,S4_OUT10r_reg,S4_OUT10i_reg,clk,rst);
Register #(.size(16)) Register_S4_11(S4_OUT11r,S4_OUT11i,S4_OUT11r_reg,S4_OUT11i_reg,clk,rst);
Register #(.size(16)) Register_S4_12(S4_OUT12r,S4_OUT12i,S4_OUT12r_reg,S4_OUT12i_reg,clk,rst);
Register #(.size(16)) Register_S4_13(S4_OUT13r,S4_OUT13i,S4_OUT13r_reg,S4_OUT13i_reg,clk,rst);
Register #(.size(16)) Register_S4_14(S4_OUT14r,S4_OUT14i,S4_OUT14r_reg,S4_OUT14i_reg,clk,rst);
Register #(.size(16)) Register_S4_15(S4_OUT15r,S4_OUT15i,S4_OUT15r_reg,S4_OUT15i_reg,clk,rst);
Register #(.size(16)) Register_S4_16(S4_OUT16r,S4_OUT16i,S4_OUT16r_reg,S4_OUT16i_reg,clk,rst);
Register #(.size(16)) Register_S4_17(S4_OUT17r,S4_OUT17i,S4_OUT17r_reg,S4_OUT17i_reg,clk,rst);
Register #(.size(16)) Register_S4_18(S4_OUT18r,S4_OUT18i,S4_OUT18r_reg,S4_OUT18i_reg,clk,rst);
Register #(.size(16)) Register_S4_19(S4_OUT19r,S4_OUT19i,S4_OUT19r_reg,S4_OUT19i_reg,clk,rst);
Register #(.size(16)) Register_S4_20(S4_OUT20r,S4_OUT20i,S4_OUT20r_reg,S4_OUT20i_reg,clk,rst);
Register #(.size(16)) Register_S4_21(S4_OUT21r,S4_OUT21i,S4_OUT21r_reg,S4_OUT21i_reg,clk,rst);
Register #(.size(16)) Register_S4_22(S4_OUT22r,S4_OUT22i,S4_OUT22r_reg,S4_OUT22i_reg,clk,rst);
Register #(.size(16)) Register_S4_23(S4_OUT23r,S4_OUT23i,S4_OUT23r_reg,S4_OUT23i_reg,clk,rst);
Register #(.size(16)) Register_S4_24(S4_OUT24r,S4_OUT24i,S4_OUT24r_reg,S4_OUT24i_reg,clk,rst);
Register #(.size(16)) Register_S4_25(S4_OUT25r,S4_OUT25i,S4_OUT25r_reg,S4_OUT25i_reg,clk,rst);
Register #(.size(16)) Register_S4_26(S4_OUT26r,S4_OUT26i,S4_OUT26r_reg,S4_OUT26i_reg,clk,rst);
Register #(.size(16)) Register_S4_27(S4_OUT27r,S4_OUT27i,S4_OUT27r_reg,S4_OUT27i_reg,clk,rst);
Register #(.size(16)) Register_S4_28(S4_OUT28r,S4_OUT28i,S4_OUT28r_reg,S4_OUT28i_reg,clk,rst);
Register #(.size(16)) Register_S4_29(S4_OUT29r,S4_OUT29i,S4_OUT29r_reg,S4_OUT29i_reg,clk,rst);
Register #(.size(16)) Register_S4_30(S4_OUT30r,S4_OUT30i,S4_OUT30r_reg,S4_OUT30i_reg,clk,rst);
Register #(.size(16)) Register_S4_31(S4_OUT31r,S4_OUT31i,S4_OUT31r_reg,S4_OUT31i_reg,clk,rst);

stage5 S5(S4_OUT0r_reg,S4_OUT0i_reg,S4_OUT1r_reg,S4_OUT1i_reg,S4_OUT2r_reg,S4_OUT2i_reg,S4_OUT3r_reg,S4_OUT3i_reg,
		  S4_OUT4r_reg,S4_OUT4i_reg,S4_OUT5r_reg,S4_OUT5i_reg,S4_OUT6r_reg,S4_OUT6i_reg,S4_OUT7r_reg,S4_OUT7i_reg,
		  S4_OUT8r_reg,S4_OUT8i_reg,S4_OUT9r_reg,S4_OUT9i_reg,S4_OUT10r_reg,S4_OUT10i_reg,S4_OUT11r_reg,S4_OUT11i_reg,
		  S4_OUT12r_reg,S4_OUT12i_reg,S4_OUT13r_reg,S4_OUT13i_reg,S4_OUT14r_reg,S4_OUT14i_reg,S4_OUT15r_reg,S4_OUT15i_reg,
		  S4_OUT16r_reg,S4_OUT16i_reg,S4_OUT17r_reg,S4_OUT17i_reg,S4_OUT18r_reg,S4_OUT18i_reg,S4_OUT19r_reg,S4_OUT19i_reg,
		  S4_OUT20r_reg,S4_OUT20i_reg,S4_OUT21r_reg,S4_OUT21i_reg,S4_OUT22r_reg,S4_OUT22i_reg,S4_OUT23r_reg,S4_OUT23i_reg,
		  S4_OUT24r_reg,S4_OUT24i_reg,S4_OUT25r_reg,S4_OUT25i_reg,S4_OUT26r_reg,S4_OUT26i_reg,S4_OUT27r_reg,S4_OUT27i_reg,
		  S4_OUT28r_reg,S4_OUT28i_reg,S4_OUT29r_reg,S4_OUT29i_reg,S4_OUT30r_reg,S4_OUT30i_reg,S4_OUT31r_reg,S4_OUT31i_reg,
		  W0r,W0i,W1r,W1i,W2r,W2i,W3r,W3i,W4r,W4i,W5r,W5i,W6r,W6i,W7r,W7i,
		  W8r,W8i,W9r,W9i,W10r,W10i,W11r,W11i,W12r,W12i,W13r,W13i,W14r,W14i,W15r,W15i,
		  S5_OUT0r,S5_OUT0i,S5_OUT1r,S5_OUT1i,S5_OUT2r,S5_OUT2i,S5_OUT3r,S5_OUT3i,S5_OUT4r,S5_OUT4i,S5_OUT5r,S5_OUT5i,
		  S5_OUT6r,S5_OUT6i,S5_OUT7r,S5_OUT7i,S5_OUT8r,S5_OUT8i,S5_OUT9r,S5_OUT9i,S5_OUT10r,S5_OUT10i,S5_OUT11r,S5_OUT11i,
		  S5_OUT12r,S5_OUT12i,S5_OUT13r,S5_OUT13i,S5_OUT14r,S5_OUT14i,S5_OUT15r,S5_OUT15i,S5_OUT16r,S5_OUT16i,S5_OUT17r,
		  S5_OUT17i,S5_OUT18r,S5_OUT18i,S5_OUT19r,S5_OUT19i,S5_OUT20r,S5_OUT20i,S5_OUT21r,S5_OUT21i,S5_OUT22r,S5_OUT22i,
		  S5_OUT23r,S5_OUT23i,S5_OUT24r,S5_OUT24i,S5_OUT25r,S5_OUT25i,S5_OUT26r,S5_OUT26i,S5_OUT27r,S5_OUT27i,S5_OUT28r,
		  S5_OUT28i,S5_OUT29r,S5_OUT29i,S5_OUT30r,S5_OUT30i,S5_OUT31r,S5_OUT31i,
		  clk_MAC,rst,count_reg,count,flag);	
		  
Register #(.size(16)) Register_S5_0(S5_OUT0r,S5_OUT0i,S5_OUT0r_reg,S5_OUT0i_reg,clk,rst);
Register #(.size(16)) Register_S5_1(S5_OUT1r,S5_OUT1i,S5_OUT1r_reg,S5_OUT1i_reg,clk,rst);
Register #(.size(16)) Register_S5_2(S5_OUT2r,S5_OUT2i,S5_OUT2r_reg,S5_OUT2i_reg,clk,rst);
Register #(.size(16)) Register_S5_3(S5_OUT3r,S5_OUT3i,S5_OUT3r_reg,S5_OUT3i_reg,clk,rst);
Register #(.size(16)) Register_S5_4(S5_OUT4r,S5_OUT4i,S5_OUT4r_reg,S5_OUT4i_reg,clk,rst);
Register #(.size(16)) Register_S5_5(S5_OUT5r,S5_OUT5i,S5_OUT5r_reg,S5_OUT5i_reg,clk,rst);
Register #(.size(16)) Register_S5_6(S5_OUT6r,S5_OUT6i,S5_OUT6r_reg,S5_OUT6i_reg,clk,rst);
Register #(.size(16)) Register_S5_7(S5_OUT7r,S5_OUT7i,S5_OUT7r_reg,S5_OUT7i_reg,clk,rst);
Register #(.size(16)) Register_S5_8(S5_OUT8r,S5_OUT8i,S5_OUT8r_reg,S5_OUT8i_reg,clk,rst);
Register #(.size(16)) Register_S5_9(S5_OUT9r,S5_OUT9i,S5_OUT9r_reg,S5_OUT9i_reg,clk,rst);
Register #(.size(16)) Register_S5_10(S5_OUT10r,S5_OUT10i,S5_OUT10r_reg,S5_OUT10i_reg,clk,rst);
Register #(.size(16)) Register_S5_11(S5_OUT11r,S5_OUT11i,S5_OUT11r_reg,S5_OUT11i_reg,clk,rst);
Register #(.size(16)) Register_S5_12(S5_OUT12r,S5_OUT12i,S5_OUT12r_reg,S5_OUT12i_reg,clk,rst);
Register #(.size(16)) Register_S5_13(S5_OUT13r,S5_OUT13i,S5_OUT13r_reg,S5_OUT13i_reg,clk,rst);
Register #(.size(16)) Register_S5_14(S5_OUT14r,S5_OUT14i,S5_OUT14r_reg,S5_OUT14i_reg,clk,rst);
Register #(.size(16)) Register_S5_15(S5_OUT15r,S5_OUT15i,S5_OUT15r_reg,S5_OUT15i_reg,clk,rst);
Register #(.size(16)) Register_S5_16(S5_OUT16r,S5_OUT16i,S5_OUT16r_reg,S5_OUT16i_reg,clk,rst);
Register #(.size(16)) Register_S5_17(S5_OUT17r,S5_OUT17i,S5_OUT17r_reg,S5_OUT17i_reg,clk,rst);
Register #(.size(16)) Register_S5_18(S5_OUT18r,S5_OUT18i,S5_OUT18r_reg,S5_OUT18i_reg,clk,rst);
Register #(.size(16)) Register_S5_19(S5_OUT19r,S5_OUT19i,S5_OUT19r_reg,S5_OUT19i_reg,clk,rst);
Register #(.size(16)) Register_S5_20(S5_OUT20r,S5_OUT20i,S5_OUT20r_reg,S5_OUT20i_reg,clk,rst);
Register #(.size(16)) Register_S5_21(S5_OUT21r,S5_OUT21i,S5_OUT21r_reg,S5_OUT21i_reg,clk,rst);
Register #(.size(16)) Register_S5_22(S5_OUT22r,S5_OUT22i,S5_OUT22r_reg,S5_OUT22i_reg,clk,rst);
Register #(.size(16)) Register_S5_23(S5_OUT23r,S5_OUT23i,S5_OUT23r_reg,S5_OUT23i_reg,clk,rst);
Register #(.size(16)) Register_S5_24(S5_OUT24r,S5_OUT24i,S5_OUT24r_reg,S5_OUT24i_reg,clk,rst);
Register #(.size(16)) Register_S5_25(S5_OUT25r,S5_OUT25i,S5_OUT25r_reg,S5_OUT25i_reg,clk,rst);
Register #(.size(16)) Register_S5_26(S5_OUT26r,S5_OUT26i,S5_OUT26r_reg,S5_OUT26i_reg,clk,rst);
Register #(.size(16)) Register_S5_27(S5_OUT27r,S5_OUT27i,S5_OUT27r_reg,S5_OUT27i_reg,clk,rst);
Register #(.size(16)) Register_S5_28(S5_OUT28r,S5_OUT28i,S5_OUT28r_reg,S5_OUT28i_reg,clk,rst);
Register #(.size(16)) Register_S5_29(S5_OUT29r,S5_OUT29i,S5_OUT29r_reg,S5_OUT29i_reg,clk,rst);
Register #(.size(16)) Register_S5_30(S5_OUT30r,S5_OUT30i,S5_OUT30r_reg,S5_OUT30i_reg,clk,rst);
Register #(.size(16)) Register_S5_31(S5_OUT31r,S5_OUT31i,S5_OUT31r_reg,S5_OUT31i_reg,clk,rst);		  
		 
endmodule
